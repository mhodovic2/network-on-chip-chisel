module noc(
  input   clock,
  input   reset
);
  initial begin end
endmodule
